module kogge_stone_adder(
    input [31:0]    i_a,
    input [31:0]    i_b,
    output [31:0]   o_sum 
);

   

endmodule
